package pkg;
	
	import uvm_pkg::*;

	`include "uvm_macros.svh"

	`include "../sv/ahb_agent/ahb_seq_item.sv"
      
	`include "../sv/ahb_agent/age_config.sv"
	
	`include "../sv/env_config.sv"

	`include "../sv/ahb_agent/ahb_driver.sv"
	`include "../sv/ahb_agent/ahb_monitor.sv"
        `include "../sv/ahb_agent/ahb_sequencer.sv"
		`include "../sv/ahb_agent/ahb_agent.sv"
		`include "../sv/ahb_agent/ahb_sequence.sv"

	//`include "reset_age_config.sv"
	`include "../sv/reset_agent/reset_sequencer.sv"
	`include "../sv/virtual_sequencer.sv"

	`include "../sv/virtual_sequence.sv"

	`include"../sv/ahb_agent/ahb_scoreboard.sv"

	`include "../sv/reset_agent/reset_driver.sv"
	`include "../sv/reset_agent/reset_agent.sv"

	`include "../sv/ahb_env.sv"
	`include "../../test/ahb_test.sv"


endpackage
